�6�   ��%�   ��5�   ��5�   ��5�   ����   ��%�   ��E�   ��5�   �x5�   �h5�   �X%�   �H5�   �85�   �(E�   �E�   ��~   ��C   ���~   ���u   ���w   ����   ��ą   ��o   ��Tw   �x�w   �h�    �X4�   �H�    �8T�   �(�~   ��u   �   ��C�   ����   �ؓ�   �ȣu   ���u   ��c�   ��C�   ��S�   �xS�   �h��   �Xs�   �H��   �8��   �(��   ���   �S�   ��R�   �肅   ����   �ؒ�   ��r�   ��r�   ��   ��   ��   �xr�   �hR�   �XB�   �HB�   �8��   �(r�   �M�   ��l�   ��L�   ��܅   ��܅   ��,�   �Xv   ��)�   ��'�   ��5�   ���   ��Ѕ   ���   ����   ���   �H*�   ��   ��V�   �xŅ   ��s�   �҅   �(��   ��>�   ���x   �Ț�   ��   ��f�   ��ą   ��B�   �Ȑ�   ��Nw   ���   �K�   ��   ��w�   ���   ��w�   ���   ���   ���   ���   �x�   �h�   �XG�   �H��   �8G�   �(�   �ׅ   �ׅ   ��օ   ��օ   ���   ��F�   ��F�   ��օ   ����   ��V�   �xv�   �h��   �X�   ��@�   �8��   �(��   �&�   �х   ��Ѕ   ���q    ���    ��Ѕ   ����   ����   ����   ����   �x��   �h��   �X��   �H0�   �80�   �(��   � �   �@�   ����   �诅   ��?�   ��O�   ���   ����   ���   ��?z    �x_�   �hoT    �X��   �Hυ   �8_�   �(υ   ��   �?�   ����   ��.�   ��ޅ   ��N�   ��.�   ��N�   ���   ��^�   �x>�   �h>�   �XN�   �HN�   �8�   �(.�   �N�   �.�   ��m�   ����    ���   ����   ��=�   ��݅   ��݅   ��-�   �x�x   �h-�   �XM�   �H�   �8}�   �(݅   ���   �8Ņ   ��d�   �hӅ   �X�   ��ԅ   ��D�   ��t�   ����   ����   �x�   �h�   ��c�   �xc�   �X��   �H�   �8T�   �(ԅ   �ԅ   �ԅ   ��Ӆ   ���   ��Ӆ   ��Ӆ   ��Ӆ   ����   ��c�   �HӅ   �聅   ��a�   �8Ӆ   �(�   ��   �Å   ��҅   ���   ���   ��r�   ��ҍ    ���   ����   ��҅   �x�   �h҅   �XR�   �Hb�   �8b�   �(�   ��   �R�   ���   ��х   ��х   ��х   ��1�   ����   ���   ����   �xх   �