{c�����C���$W� �D�m-���b5���
V��&~)޻��EdO߀y�V��3^���k!����5a)@��\�vGisat�!��t���6�R�	�m��+�^v�Y?:�0/�]U�	uj�L�ä��@��`y���ٝ�ʁ	l���5�L3��Y�;�jXx�d�=�\�b) 1�0�ƃ��;zD����m]e��-�m3����A��ic�    �#���]%ͩ%��kի|SG_ʥ�O���ć8��c*��{��RC!#�� ����<    �&Lu�E�I!ߪ�����8�WI�jv �wQ�$�!�M"�%ݍ���Px�Iʆm    o�*|ɃY�h�ZR�J���h*�y��&:W�g�?�̩W�,�����9"����aE��g    _�L^��
\u6w�
�a{΍���lO��l�x��W� Db��-��bL���q˰^��)!    OZ	ܵ�S���bkL�p�S�oa�̇��~�GD0�t�D\�ͨl����"��W��I�    ?u�N$�U�MjQK[&�R�>� я�z6E#7�,�R$_X}"£@G�w����	h�u    /,"I<R]��{2�钇K\�`(V�A�6�|f['r�$Ԭ�M}^��r����	�V@��dye�_�B��|�l·5�z�̇�;�s�X���J�뽗3���e���q"+e��{p;����`n�NwnI_��f�@�z�0+�8��e!B�VFf��g04%./]�3 Ҡ㣥Z�`"Y�g�U)��gP��\>��)*x��&ͩ���!��u��:x���dC?��YТ��O�=�1_�ŕ�Τ~�w��M���+��?d�̿��jW�e;��ց����M��=PxM2��0��� ��u9��B~�C����:,��O�I./�S����_}^��q��pV���N���CHӭ�(��K_s�10�g���5C.����A��\G��e�fO:�� �+�[H}B�w+���Ǜ/��%�-�^�o>lc-�y`��Bb���OY�<���?<z��K�^d���Yx�3}Q�� �q$��ۮB�QS5���.$������L���/���E/ �Vʑ���Ψ?f��zޛfBg���T��������"C��[ǰ��V�>8Rҟ��s� �s�2J�5��m���|�1�Z1;8�*_��TI�md!�(O�3�a�4IWi��Y�,�
�����$Q%���)�׫;���ڕ�m�*�뷒��I#��l��B�R�6m#uS� �K��/�o��"�@��LX�ѕ�.�����e �8��#[�v�8[w����dqM�]��W��sP�Q�I�swN��(oG�|lr�)��Z-����!�hԷR�Pm�&�ؐg����i1�s���|�A�g�Ȟ���-�R�8_���gGu]d�
���{�H�'���[*��r�W�yD%)�-�w�bG/��p���Q5)����w>}O)��ؕ^���`��k�uȦa#��Ρ_G�u�tgB�����M���|�=��ذ�݉v^(��?��1�hU��jl�[�s�Q��Ѧ 16��&7<�C������.��dCh~	_�eC]/{P�<�&.��m�T�K��()�A�P��'�^�ԯ��}�KPr�O��(��@�Hyrɾ-�H�\�l%�H5���g� ;�ŬX,0U�