c a l l ( b , " i n t l " , g , { h a s h : { } } ) : g = h , f + = n ( g ) + ' < / e m >   < / a >   < / l i > \ n                         < l i >   < a   h r e f = " h t t p : / / w w w . a b i n e . c o m / p r o d u c t s / m a s k m e / s u p p o r t / f a q . p h p # w h a t i t s t o r e s "   t a r g e t = " _ b l a n k " >   < e m > ' , g = " m m _ h e l p _ w h a t D o e s " , i = c . i n t l , h = i | | A B I N E M A S K M E . D u c k b o n e . H a n d l e b a r s . g e t A t t r ( b , " i n t l " ) , t y p e o f   h = = = k ? g = h . c a l l ( b , g , { h a s h : { } } ) : h = = = m ? g = l . c a l l ( b , " i n t l " , g , { h a s h : { } } ) : g = h ; i f ( g | | g = = = 0 ) f + = g ; r e t u r n   f + = ' < / e m >   < / a >   < / l i > \ n                         < l i >   < a   h r e f = " h t t p : / / w w w . a b i n e . c o m / p r o d u c t s / m a s k m e / s u p p o r t / f a q . p h p # l o c k i n g "   t a r g e t = " _ b l a n k " >   < e m > ' , g = " m m _ h e l p _ h o w P r e v e n t " , i = c . i n t l , h = i | | A B I N E M A S K M E . D u c k b o n e . H a n d l e b a r s . g e t A t t r ( b , " i n t l " ) , t y p e o f   h = = = k ? g = h . c a l l ( b , g , { h a s h : { } } ) : h = = = m ? g = l . c a l l ( b , " i n t l " , g , { h a s h : { } } ) : g = h , f + = n ( g ) + ' < / e m >   < / a >   < / l i > \ n                         < l i >   < a   h r e f = " h t t p : / / w w w . a b i n e . c o m / p r o d u c t s / m a s k m e / s u p p o r t / f a q . p h p # t e l l n o t s t o r e "   t a r g e t = " _ b l a n k " >   < e m > ' , g = " m m _ h e l p _ c a n T e l l " , i = c . i n t l , h = i | | A B I N E M A S K M E . D u c k b o n e . H a n d l e b a r s . g e t A t t r ( b , " i n t l " ) , t y p e o f   h = = = k ? g = h . c a l l ( b , g , { h a s h : { } } ) : h = = = m ? g = l . c a l l ( b , " i n t l " , g , { h a s h : { } } ) : g = h , f + = n ( g ) + ' < / e m >   < / a >   < / l i > \ n                         < l i >   < a   h r e f = " h 